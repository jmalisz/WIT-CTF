BZh91AY&SY���� v߀Px����߰����Pxz;�v�gwvw��%F�0j{I6��0�MF�� ��?AG��F�Q� z�   �
#D�ɓ�C54 �4�G���Ph �@4� 	$j15&�6M��O)�OS�P ���(�q!(IX�\�O���(]��o�(;�ZLhM�{!�ӂ ��,h�p�jb-h��kV�����h�q�O��gDUG��6�%����m5�0���1��P*���o¡X��@�EI�i-¸S��gX@���ɇQj/L{��!��<��-�b�-����ބ��b�"	a>6]�L��<FERot̛Ha�����4�9��k.ka-ͼ:JKx��ؼi��6�l���^b��?1�Z��JΘRܲ�tv]~s�Rd14�d��1��<(�m+SE�m��{I32�g:��,���Ϥ�J<�M����'u?V4M��u
`P��F���Ft�Y��*OB�9ب�����8����M�2�Pj/�u�b�)L�+Idאp��]�D�0�/@�y7�f�&\Q����R���OM՘bQ.h��'AS\�2�XYP5TQ����uM�g"!��kͺ�,P���d�i���bF[}J�N#�I�nf ���gTL�TҤ4�$Z�)�Zo��F�Gv���A"�k��BcH�:̸��WWR�jS��[9_s��QJ
5��bVR�$w��Ýpl�%n΂�(#�)�D(V�13�̋�l�S�<Ӳs�N��!)d1��^�QܦGI3T� cx�I�ZLA�=��AB2�,/b� �=tNl""A(3����
�T�K�a�")��ni�6���x�^�Q�A ��E��
)��!�2+�l�%}�<d�I���N�7"
�bv��8h$OE�஬*x&q��1�b��R�+����\�UD�+��ei-	���l~�E��;N.rE����"���%I�V��`�f]Ǳ�����X�FYk��2()�h�ֻFt��#U�����g�4��=�zX"��,T�d��?�"��h��II���Jl�(J+���l\�g[^0�� ��Y�K�uX��ܑN$-��-�