BZh91AY&SYƴ7� {߀Px����߰����PxG;�v�m�uݮE�M��h�=��d4�4� &B�=G�d�4�hM ��F��&(�ѩ�	�  11�2b`b0#L1&L0I#HҞBz)�&�P~� �z�G�J����5��;.��ݑ��ޘU�Ƅ�2]vA b�9�4U1h��kf����/��}Jz��&xb���9xq.+ň�k����7v��ƴB�f���ܛcHW0x��p�b'Wy�,Eh"���n�������QT`��pnÇ��r�T��Ŭ^�1���T16C�3��D�Pi�kK
3��#��V�D�1Xs�XI�8��<����f��7��̳���@�m��r��}�U�i종3�
[�PwӶ�-J�K!P^���+0ǎ!ڄiY4Y����3!�\�������Q��ŢMg�5Oј~�򚡥��$��^���S/��3�3�icÀ[tgҎ�:�J����]&1ܚ5�	�=d5*T�����k�:�0�6P3A_��g�t\����USO����1�KI�����p�7�^e]c.H�@��#���q�}[$D8Ms��y�L
�{�@�D��*�2R� p9�c���!��
,�!LεF�Ӧ�U8S<|XT��,Q��X��C�ۦli����ť!lWu� �Q4�21C�X�Ǒ�]���w��pƥJ�Yu7������*7]�4�]|s
��G"�[��-F��Y3��+Dŕ�y;F�/�zƳ��W�����YP1��=vS� qQ��tYH��	�bt_��qT���ހ���ة���q�"(�����0����娉�0!�E�0 �^92�Q�H�.wyI�6m�`�(�C �Z�:"kˈp�R��}��ժ�	�u0�'��`%e�%��a���X�4�`d��̂�0�u���喁�6�հ�A	�uoe��󻟆4�ԍ6a��R;m�?j2h�"�V�P��e��E*AqiM�u�DT�0C=M$*?�K�Pa0�*L�6	7c4�"�y��aR/��
u��*CSN0�:�P��:
d�W�.�p�!�ho|