BZh91AY&SYSp98 �_�Py����߰����`^�$�@T�*Ts F	�0M`�Ls F	�0M`�Ls F	�0M`�Ls F	�0M`�L"�@%?Hڦ�j4�dOI���A�m#�� HОD�x�S��$ M4=A1�q������I���C�؃ ����{Zh�A,! $"9�)�{������1q��X������+��e^��Nл�6�8��t��j�+���Zw_I�Lv�6���!�{!,�M[vhfG^��	��@`Ď�fҦf.1�H��)�G%��@���@P�or6����|�y�`�1E�;������Q|����m��{��+XQ�3�V��E0�U����bSi���&�M�ɢ��d�0׬�D�0����iS����:$Q� �H��fc�424�5�.������0{�N����I#$�DK��xf��L�XS���ه��PX�kAb��+���=021*��2#x���0 ��M.PB	�����d�v�8:QA�x���X{��я�~Á!�d�3-���~�����>5���3{Q���ѹtou��T�����x�߭���ɨ��6�ē�|ߋ���2�P�`��������z��p}z2f���ݑ��C���������&�b!���=aOb����:0y�ٻ�v�$�H���a�.}�̦�?�ۆ�Z��'!&�
�swG{����f?W}���8��w6��%̡�A�7t�l,�ȅ�| �lqw��b*�p7;�(]�.v�\h	~�B4��w98�	��jG�ܖx� I�Q�y�M �h=��8bmwr�Ź�d�����>1��H�t �8ld����8�ҝ^��L�.�C��(܍�3E5�^��`Z� M�^y:Uh��У�t����gۑn���;���y��s;r(��у��ܴ A4��f�8\��̀\�� \Bn~c�Qe�),���ME*�͘�{jp3 �5.�k T$vC��F+���R�.�dp�9�����+7)^��{�������D�0u5��j'���g�A��TN�$��m0kfI�Q����[�����Q�l/C�s�rU�ͅ��Q0����`�'�q�mSj`8�`u�G	p�炷�& �湱�V����Q��a7;�P7��ŵ$��yid�Ǚ���jh�&,��-L�7[����ͩ���� �&b�)�ta�&<o�� ��Ҙ48{�n��|�dh���hn	��"�<�a�����!:JG��N��@�9�����]��BAM���