BZh91AY&SY��FB �_�Py����߰���� � �����j�	Eq�&LF& L�&@F ��Tdh h       q�&LF& L�&@F ���2b10d�2 h�00�L��O55='�ze=�h�4��4�$!CT�ҞH𧩰��P zF�4��E(C
b���l�|ܑl�w����Au}�Ȑ�b,BhƘ��l
7��=��2��B�G��OZ���Qj��>�u���|���I0��u��9�%;�
=�f6`:����8��֚�d�%���߮�{�"#'4$��۲���[o�]ZԼ���)\�(b���4�e4Eҍ�Y,��t�)s�^�|���LaeF�b��.�4�s��d����5;ڍ�i�s��b wζ�r�[a���͒0��M�%�Vo����g`�b4��n�}�tWN��HM6ٲ_c:Ni�Q�,�a��vf���t�;�=��w�$0h�w�K���+N����{l�SB!��2.������
��v���HB2&��P���BL �0r����&�ϲ�l0ӫ���=��C��'��BL�7�I�)I��qC6�{$-(\��������AF�6��mB�I����o�)�VH���g�ڒ%�ve�W#����D�h�C'��b'��P�P�_�L�+�x�t?$(<���?�[��=�4:�}O#Ƈ��C��N���C iG��c�(u�=��&�i�f��v�n�c]3�C���޳��ڃE��?'��X|�+$:�!40x �f��@B�K6�2|�u���AV�~o`M��	*I�X�{�����P�ס���u$6>t-���D��z�Cv:�$H��6V�L8rz�>��u!�@�!3�K���D4�⛟4��x���� B!N(b��>0y��C^�A�u�D�rp��֏��|�� �C��
�C7y�P��\��Ws]���ЇpS�9��7B��tN�{�sa!I��4�CR(w�͆����)a7i���P�c�H�DiC&X�Sd�ץ��d��^M�L׼�ݱЇ`�Z)�nTd}7Ѕ���HI���6��'f!HSw�������,;�{ڇ����ӡV�h�qQ�F!VN��}���慃h>Q*ڎ�֨�q�B� ���[V��
2�s0Xk̉�o6�Hg��2<ܛ���t	�6��96.hP������<$���Q�sG`��|m�!D�y�HɅ��
^�A}���p<L�օ����d=q"�]�(s!;^@}-�H8���L�ܝ��?��7����)��r2