BZh91AY&SY��α v߀Px����߰����P}ǧ�y۷R���$�I�2OOSj� A�4 R4��	�3P CF�@�$D#STh�ML�OP�=F� � ��j=&�6��� hi�   �!4Ё6�Q�x�d����']h�V�hY�A�@�}�.�9Nl�I�	�1d4�.� .�h�h�b,уR�wg3��a�>U)�:d���h��m�W+�F���a�z��Ƹa@��G��o�����@p�R8d��:E`���\`Y�����f�%Q�c����{��%��&�wQS=+��ĵ�,��,H�^�x�Ͳ��35)�D!M���gRd��mZ读��ʨM���ܳ�����d'b��{�Y��颅3�
[�PxS�oK5������(5�Wa�lC���4]���o��Z�1�UeD�e<5��0+�v-����h�j��:��O"�Nڠ���� �7���D�.�o<�i^��i#%2b���-Ǆ���j��ŀ2E�_�FtD���U��.�e�K!�@�q����=V,�2�s��f����^9 r�
`UDG(���� '7( ����I	h'�R�d~ɳ8a2��eۍ�8ʨS3�Q�D4�Y<�T�͔�X,V���!i��<]	��芹sA0��e��u^R�d[ho�zP0L�8�
Է�ly�7��I s�i	�=�A��E��h���:Y1�ƌA��jO�N_fD0���Cg��8��6�ʵm��]��t�5��Ό�� ��Uf�:.��[
,
�E��!����T	�B�e2Qs��ȏT����Cmgpn���.�+@lU�8�`���j�p;�%B���=E��2*1��QK ؐ`D�UXD��̐u���ׅ8-z��:������T�uwM2)!�ۨi'����+b́�PX3���w3�:J,�,;��X�RLlӊ2�6�H�	�9u�Y�C�LtJj���Pr�M�.C�[䷪��G�FK	J�$`����#k��Լ�f�K�9y\W��Eь��z̝�Ʉ��Ԧ�ϛcm������K21H��rE8P���α