BZh91AY&SY��Ã ߀Px����߰����P�����v%�IM5457��D�M�2 �i��@���iL�zM�zM4i�� D��z���Oj�Q�iQ� ��d0	����L&i��H��5L4�I�i���@   ��X
PJİ��D�8�����p�T`6+\4p�P�sF��TiU����_�nȅ�62y�D=~�.���BL���*x9�`p������m±�$��(�;�J�@fZ�������cѳT8w��ib�h���~��Tw�s(����q���;e��h�+�F�&�Tb�'�D�pa�"$[~�k��K�vt�cO���Rڹ�[�"��q>3 �����*�v�j��P���\�ca4Սc���+�fݡΖ�rY`�}F�����(�Q�$^�%0���C1S������]�c�K);Ơ�U��Jrj��c� �~j���`���j3�f��S�U2yg�O�~��[
�eut���c��odf�S(���0����0���f��~h�lJIe��	H$���!�A�Ҝ�+2aj��a���\�?�~RWk7)f+�@�l�D�D~hSjA�z�eɍX��������d����xG�=6�1k�JL�a9r��y�ʫ#M�����8�lzU�w L@R�C[���	E$T<��P�d�-�mu`�Z+ņ.!��H��L�Wƙ�
)4��ةR�Mm�繴ʊ�O�)����]�JBs�1�1ezMy$����
E�1
\�Eǉ4q��6���@L�X/
����S�D��S�`-3�L3�0�1�^3���T��Ӵcgj�)!U�2/��D��E-���Z���8����;�y�0ڬ���j%e[2����5������a��6=+�y5��0R����qH�誂�#Tul��0���<X�>�bad��q	�*i���]��BC�