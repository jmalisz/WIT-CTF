BZh91AY&SY�A& p_�Px����߰����PV=(�v�rݺ��H��jM��Si�� i��  hJhК�C&OMS#j�z���A�z�	�Py�SjmM�6�� &@4d���`F�b0L�`�&��?RmO$�����6��h   �|5!&I:AD;�>�$��Ê��~�pI�	�1d4�n� .�h��Ɉ�FK[{�O�ل@2_
���RL�R;��[;�Krd)�k�0�z�Ʒ�ʑZ�͞o�!U��P�K�fFx���*	�@��prĭ͟���eQ�c�ť�C�xج��j����i�\n�bo�r����s���df�������pr�cI�U*I^�"yY#$F���;i��� a<�X?���"��H�U)����e�:��ޖ�����T�M13�0.�/C�M�dы]����X�vyN��Ɠ�R�����WH�����>���S�s�#��ba�S.����k�VQ�t$�1��;~| �	��\��
���{��=�
r�!��~���$!�Y��|��"��9�iU,h���V@�K/Q�1���^��2�T���)�*�GT+{��Uz�J��e��E/�U4�a��x.�s���& ySjhT�6�4�4Y8S;x�\��o	P������Lh�.�AL��s"�iռkbw��|� `��p7�%�1�g��@1���%^[J�r�����%�*uFVL[w{h�6����9���阆9��c(�,X�(����+1�Fkl��q_]�P���aC��; ��ӎID	���W%2Qy*g�I��pi�6և�a4U2(���O�4j�6Y<of.J�J�	4��Ό�o���6t*t�#�X�$bd�Y���cZ�L�Tߨ��Yq�$�C �#f�
�>��+ 6�d�Ap�/�i�5i+.:����+�*M(�1�w��<9Y@Տ:1ǟ!A�W�$��(F��.�4�25#��;�eU��d��P�P0>ɵHU��ޝ�%�2V��%�]��+#��˥s&F�
\	� �ͤ0�n��dB�H)��W���)��	0