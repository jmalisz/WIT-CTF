BZh91AY&SYW?�) A߀Py����߰����`_      `�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L��`�1 �&	�!��L����)��i=x���SM4���� ��L�}��}��͑��ˑ_�e��Td�R��)H�E���Ԗ��I&*G�,�2��*��.�������k3�]zz���r��`�gog
�}F/kT�I��)v.ޚS�ҕixrr�̦�*��LT�����b�ll��0b����{ �Y� �S�.z~O�v��e%UW+��YK)�}J]Q�N^g��r�r�l�s�Ş�3^SֳK)Yiu6S����G�����-{�l����|,��Q�Sk$���9��1�L����1_�nߋ|i�ne���ݏq<'B�*W������0z��h>e4}%�)��f̈́�����ԥ�`��?L�5��*J`�K,��]�s�?b��&ǵe�Ղ�U�Z��Wr��������/|���ώ�_�k�����1}�Y?�|�2����.�blX�9��M�E>/����-�6��ئ	vf)g��?��X쌖9��)�=�[�M��~�^�]�'�~1���Ã��;I�4F��9	T�x�e�l��֛�O���G:��aw�NG3�<eK�$|視�N�qW����Rx�%���v�H��x��1MW<�$�I�������h8+,�CM�SIjV�p��.ɒ���������Yܩ.��\����]u��C���2���3��j͡,c2����m)&Y���z'g2Q��N,f��d�M��OI��dͪY:F���jw�ϻ�˻
��%'*�e�a��܏P����S��֘�yS�`h����E4I��Ι�R�t�8��j��k��'��Y��O�p�}���z�fЧ�����P��sgi"��$��V�ک8J.���Z=�dng#]�)#j`���,L96*ʵ�KKúģq��-��'׉ʺLOqvs(Z���R���%�CX�3�-�޹1�t�WO����j\����/#@�ށ��b^O�RJo��Xqw��3�l1O��Y�>,b�I�E�,Z`�s:�'\�mT��ΉR�����hb�J�Sz���T��$�S���N�Q���M������4��$���iI�ѣ&X>�1WB�K�s������fY���5LOɛ/��'2nM��C3��u��7,n;�p��6m��	�g"���c_���rE�.�D�609$O���&���Xr����uKG^3���:#�`��)�R����x.Z�t4m���.�p� �R