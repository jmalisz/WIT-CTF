BZh91AY&SY���[ i߀Px����߰����P}���k�Fm���	"C �����z�M��h �C�4�$�U?Bi4�d�� &!�0$D&P�LL�i�3S	�  i����L�L�@d@    �Q�~@��mLdM<����  ���E�iP�|�ԋ/����퀳	1�6�.� �1Z9�4Y1hɩk�{K�6e�9R��$Ψ�#����Kk�cT��skټ�5�
R�����V�X�4)�J�Q\V�� Z�X4�~���YLy�����9ܴY#���36Ѵɇ�n.T4������
��.�z�AW0�	��-���#�o�ţY��ǥ/�m��	�\b�?���"�䰫5쪅3��,���׊𫈅h�
)2lgh����(@6��F�v�ڻXgA����Ym㢿⸪r��џ��aγ�Ѯ�N�r�(�ۚ��n��D%E�����������:�Y�b�Yi�<(��]��z�Xe�9��#���ί�`��2��+;���;���a�l��Kn1<�.lq�70)�jᢾ�F��(����:\R�h�+�|�K��Z$f@��,#��!:�$g���UTCN����j��������s�!�EH�&2�銅}ˈ�� ��b����ҝh�HSt/B�����g��8s��̋��j�*Ӂ��X8�O���dv
�!��g�Ɋ]ޔd���\Ṫ<�mr!�rJ2�eRի!a��I��t�cY(��Jb+��'E�2aL��tz���j�t�A��P��L�]56�Fr�E�M�a���尉�0�+@p��Ȋ���ٔN��	HKv:��fR6aF�R��&��8�3I�q$�}֧�r��L㩱r܋��-"�:j��!1lZ�+(�[p�&!	w������1aJoJ�0g�
X
A`~I���20뀠���&�b�xq��u�?�T����&4`V���T`y�Z�&�\T"��u��Q��^�u�6W.�����ѡ)�Tܾ�e0���^d��	����(d�d�J��$��w$S�	.��