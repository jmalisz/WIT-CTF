BZh91AY&SY�Ú u_�Px����߰����PV��wS�����H���M��Lb4ѡ� d $�m$ڧ��=�&��ɧ��@�	��I��cSF�=M3Q� @4d���`F�b0L�`���������S$4��   4T�vhI�P�Q/���N��r7�~��&4&������ 1b�9�4Y1h��k����M����mJ}��$͢�;Z���.-�!H�ֿ�n�jc�u�p���s�i:�t��j�G0�� E��o�"�k���e��0Ly�pÇ�7L
�s��Y7�&t�<4���bl��Y��0���s`�شt��I��������
1��F�զ��,���&u���Z�Op�m�ƻ僨{�Y��Wޔ)�p��e�+�~5{�PZB�&�E�X��lC1�iY4^�X���b���UR|�)���~��.��N:��_Q����Z�Ɇ4k�I�|;(��vV4�S g_ˋE�7Z��&0$2��Q���z���i�v�C�Ј�R1�.�	�\���ն5���wVQ�D�՚C
O��k��pb)ł��K��S��]��$��4FTE/�V�I��|C/a��>l��ǕlLUOpE!�Yœ�9��f7�q��y�ԏ���n2aL,�W

�=�*	�yS��
��Cyv>�*?FI��8dS���ϽU�*& i����&��R@Ds��JV�EXT�d���2/��R|D�2�F�T���!�Z�1�V����LԬ���I�m� ⢼��N��++afC��P�/L���gN9R�&o!]��)t\h����oi�6֗�a4V�Tpܣ��2΋!r��=�[�v�1D�[���Of �$)v$q�QYK��d�,�ubTA3��F��%�|��
K!pa�lט�+��Y�4�C�z�ѫ��a�X�hx��YX�4�'��L�\���5�r.-��e ��L^�=���&b1�P�]�yͮhPk';&�0>����ZS��˕:V��%Ѿ�i��kF��tw!C&�5(��=��o:�(�=��-�{�]��BBYW6