BZh91AY&SYBqt� x_�Px����߰����P{�]6sn�KM:0�H��6��6��ȍ���dh  4�&����=M�hh�4�A�D"�
z�(`�S����101��&$Jh�DMO��č��  �J=��JVH1 ���a([9�DPv�i1�6���ֈ �A[G&"�����8_ѳ@j)ʔ��Lꊨ��ϫ��%�H�#]�m�q�kM�H���<ᎡY��%M��k��@̼%����]LE��1�ٙ�C�8�P&�[P�.n�˜q�J�!��B��4�"�3|22G�&��P&pS5J�%�RB�( �K-a�6����Ci�� a>�.���"��Q[)B��-�(x@���6���`�~�]�!�"iQ4Q�g���@�&/:�׺����}PQ�S�-nϔ~��
ƖآL}6I�|�^�(0��Bk��˳��k �L�0���,G���:+�=�T�u���:�(}�V�`�*e�@�9�\3�X���)�Z1�K��=�5v�ʃ�H��A��UF
��C$jh1���X# �5[A�� LBe��e��:ldݎ��J�M
���4�,]8UU�l�&e���
��26s�f#S�T��`_u$��[I
Ȇ��ޗ���H� �ޯKr:eڹ3�Rpz�DҳfҴ��UlX�)EJ�C;&&s�21�~�^���z�B+$�,JAc�X��	\�fʭ@��l�֔ʠXYi�(F)���I��RG��Pp��Pp�����)����zDRN����X>�E��B&�ҫ�	��.UՊ �Tۭb��(���G ����0"���h�XFL�b0�H��E��U+��8r����ֹK��Iu4tn�S%�(����]��p/���5�,(u�Y�\7�R�N��Y�ˁU/5=V��q��T���C���l�K�uau�D�f�{��U���裭
��N
�[T%t�]��+�Ў�bǡiP�U��b]�u\�J���}0����D!bȃ=����ܑN$�]0 