BZh91AY&SY�N �_�Py����߰����P�ye�	���Jzi��ji�SML����4z�h1�`�1 �&	�!��L�����i2���M��ꌏ(4  G�`�1 �&	�!��L���#&�&S�S4�F��f���Fh4Ԕ{�A%	*�,#���MRP�z��<P7&0bM�{!���D 0iZ<.M"�5-sqr���h�v�9R���*g�)H��z'!���R5���5��l��n��EG�z�T05��"�aC���bw!���hKJ��
��"����f�wv�;XQ�[��1b�+|�w#���d��m��2ŭ�A��q;�z�P��(�O���<��i�<�Mq��M3y����pƁʮ�����1���m��@�+�w�"��U���B��
[�P�������HUI�n3s�;�BlFo�����4�fmwAkpa����,���Pq�����p�Jm~�K+Ȧ�G�Y��o����:B9WC�	���||Z�f`�)�LwG�y�*9O*�rx]����uY�`v����CCi* �i���S ���n8.(�tuN�Q%^n�E��7�P�ڋ@5'L�S3���a���6Q����m��B��]VE��^Ec,��*/i詛Tq�K#$�&u�Js�\�)��mq`*`�#vA8�"��%|�X&4
�?�C%^m<E�0�I�=$�F�؆>�|��@�s�8�d�����RT�Cd%jZT������!���0�2b�w�Õ]�=W�s�^��ḪF�!����,ucS�31�\1��Se�b,#3��=��銌KQm�T��a	A�	�ʤ��L�^*��D�K��0���}�e�&ȘTA�pܩ�y$�V���4�oG?a M�Z6�A� kq,:#�-+�\R�I���j[�8��c�~K��-e��jdm�`�Q0��pfa��qy~�^DJΒaX�Ç� �B�D80Gg%��iO���:Qv�ܨ9פ-'1��k��2���9"�1�Ý˂�".FqZ���&�J9�\��[�������b���yoҝ�T�a/���L*��a����3��Y���;��ܑN$�CӀ